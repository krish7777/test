`timescale 1ns/1ns

`include "mips_core.v"

module mips_testbench;

	reg clock;
	wire result;
	
	mips_core test(clock);

	initial clock = 0;

	initial begin 

		$dumpfile("mips_testbench.vcd");
        $dumpvars(0, mips_testbench);
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
		#100 clock=~clock; #100 clock=~clock;
end

endmodule